module mux4_to_l (out, i0, i1, i2,i3, sl, s0);
output out; 
input i0, i1, i2, i3;
input sl, s0; 
//??????????????? reg out; 

endmodule